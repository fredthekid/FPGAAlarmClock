module timer(
        );
