module display(
		input wire clk,          // main clk
		output reg an0,          // enabling and disabling 7seg
		output reg an1,          // enabling and disabling 7seg
		output reg an2,          // enabling and disabling 7seg
		output reg an3,          // enabling and disabling 7seg
		output reg an4,          // enabling and disabling 7seg
		output reg an5,          // enabling and disabling 7seg
		output reg an6,          // enabling and disabling 7seg
		output reg an7,          // enabling and disabling 7seg
		output reg ca,           // lighting up segments for 7seg
		output reg cb,           // lighting up segments for 7seg
		output reg cc,	         // lighting up segments for 7seg
		output reg cd,	         // lighting up segments for 7seg
		output reg ce,	         // lighting up segments for 7seg
		output reg cf,	         // lighting up segments for 7seg
		output reg cg,	         // lighting up segments for 7seg
		);
