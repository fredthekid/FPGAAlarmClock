module speaker(
        input wire clk,         // main clk
        output wire speaker,    // used for outputting speaker
        output wire vcc         // powering the output
        );
        
